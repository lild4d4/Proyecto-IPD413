** Voltage divisor **
.param vdivin=3.3
.param vdivout=1.2
.param vdivratio=vdivin/vdivout-1
.param vdivr1=1k
.param vdivr2=vdivr1/vdivratio

** Load parameters **
.param loadr=36k
.param loadi=1n
.param loadc=1p

** Amplifier Parameters **
.include ota-parameters.spice

** Bandgap Reference **
.include bgr-parameters.spice
