magic
tech gf180mcuC
magscale 1 10
timestamp 1691437249
<< error_p >>
rect -658 -6480 -644 -2920
rect -580 -6480 -566 -2920
rect -502 -6480 -488 -2920
rect -424 -6480 -410 -2920
rect -346 -6480 -332 -2920
rect -268 -6480 -254 -2920
rect -190 -6480 -176 -2920
rect -112 -6480 -98 -2920
rect -34 -6480 -20 -2920
rect 44 -6480 58 -2920
rect 122 -6480 136 -2920
rect 200 -6480 214 -2920
rect 278 -6480 292 -2920
rect 356 -6480 370 -2920
rect 434 -6480 448 -2920
rect 512 -6480 526 -2920
rect 590 -6480 604 -2920
rect 668 -6480 682 -2920
rect 746 -6480 760 -2920
rect 824 -6480 838 -2920
rect 902 -6480 916 -2920
rect 980 -6480 994 -2920
rect 1058 -6480 1072 -2920
rect 1136 -6480 1150 -2920
rect 1214 -6480 1228 -2920
rect 1292 -6480 1306 -2920
rect 1370 -6480 1384 -2920
rect 1448 -6480 1462 -2920
rect 1526 -6480 1540 -2920
rect 1604 -6480 1618 -2920
rect 1682 -6480 1696 -2920
rect 1760 -6480 1774 -2920
rect 1838 -6480 1852 -2920
rect 1916 -6480 1930 -2920
rect 1994 -6480 2008 -2920
rect 2072 -6480 2086 -2920
rect 2150 -6480 2164 -2920
rect 2228 -6480 2242 -2920
rect 2306 -6480 2320 -2920
rect 2384 -6480 2398 -2920
rect 2462 -6480 2476 -2920
rect 2540 -6480 2554 -2920
rect 2618 -6480 2632 -2920
rect 2696 -6480 2710 -2920
rect 2774 -6480 2788 -2920
rect 2852 -6480 2866 -2920
rect 2930 -6480 2944 -2920
rect 3008 -6480 3022 -2920
rect 3086 -6480 3100 -2920
rect 3164 -6480 3178 -2920
rect 3242 -6480 3256 -2920
rect 3320 -6480 3334 -2920
rect 3398 -6480 3412 -2920
rect 3476 -6480 3490 -2920
rect 3554 -6480 3568 -2920
rect 3632 -6480 3646 -2920
rect 3710 -6480 3724 -2920
rect 3788 -6480 3802 -2920
rect 3866 -6480 3880 -2920
rect 3944 -6480 3958 -2920
rect 4022 -6480 4036 -2920
rect 4100 -6480 4114 -2920
rect 4178 -6480 4192 -2920
rect 4256 -6480 4270 -2920
rect 4334 -6480 4348 -2920
rect 4412 -6480 4426 -2920
rect 4490 -6480 4504 -2920
rect 4568 -6480 4582 -2920
rect 4646 -6480 4660 -2920
rect 4724 -6480 4738 -2920
rect 4802 -6480 4816 -2920
rect 4880 -6480 4894 -2920
rect 4958 -6480 4972 -2920
rect 5036 -6480 5050 -2920
rect 5114 -6480 5128 -2920
rect 5192 -6480 5206 -2920
rect 5270 -6480 5284 -2920
rect 5348 -6480 5362 -2920
rect 5426 -6480 5440 -2920
rect 5504 -6480 5518 -2920
rect 5582 -6480 5596 -2920
rect 5660 -6480 5674 -2920
rect 5738 -6480 5752 -2920
rect 5816 -6480 5830 -2920
rect 5894 -6480 5908 -2920
rect 5972 -6480 5986 -2920
rect 6050 -6480 6064 -2920
rect 6128 -6480 6142 -2920
rect 6206 -6480 6220 -2920
rect 6284 -6480 6298 -2920
rect 6362 -6480 6376 -2920
rect 6440 -6480 6454 -2920
rect 6518 -6480 6532 -2920
rect 6596 -6480 6610 -2920
rect 6674 -6480 6688 -2920
rect 6752 -6480 6766 -2920
rect 6830 -6480 6844 -2920
rect 6908 -6480 6922 -2920
rect 6986 -6480 7000 -2920
rect 7064 -6480 7078 -2920
rect 7142 -6480 7156 -2920
rect 7220 -6480 7234 -2920
rect 7298 -6480 7312 -2920
rect 7376 -6480 7390 -2920
rect 7454 -6480 7468 -2920
rect 7532 -6480 7546 -2920
rect 7610 -6480 7624 -2920
rect 7688 -6480 7702 -2920
rect 7766 -6480 7780 -2920
rect 7844 -6480 7858 -2920
rect 7922 -6480 7936 -2920
rect 8000 -6480 8014 -2920
rect 8078 -6480 8092 -2920
rect 8156 -6480 8170 -2920
rect 8234 -6480 8248 -2920
rect 8312 -6480 8326 -2920
rect 8390 -6480 8404 -2920
rect 8468 -6480 8482 -2920
rect 8546 -6480 8560 -2920
rect 8624 -6480 8638 -2920
rect 8702 -6480 8716 -2920
rect 8780 -6480 8794 -2920
rect 8858 -6480 8872 -2920
rect 8936 -6480 8950 -2920
rect 9014 -6480 9028 -2920
rect 9092 -6480 9106 -2920
rect 9170 -6480 9184 -2920
rect 9248 -6480 9262 -2920
rect 9326 -6480 9340 -2920
rect 9404 -6480 9418 -2920
rect 9482 -6480 9496 -2920
rect 9560 -6480 9574 -2920
rect 9638 -6480 9652 -2920
rect 9716 -6480 9730 -2920
rect 9794 -6480 9808 -2920
rect 9872 -6480 9886 -2920
<< error_s >>
rect 1792 4071 1803 4117
rect 1976 4071 1987 4117
rect 2160 4071 2171 4117
rect 2344 4071 2355 4117
rect 2528 4071 2539 4117
rect 2712 4071 2723 4117
rect 1792 1959 1803 2005
rect 1976 1959 1987 2005
rect 2160 1959 2171 2005
rect 2344 1959 2355 2005
rect 2528 1959 2539 2005
rect 2712 1959 2723 2005
rect 306 1521 317 1567
rect 363 1521 374 1532
rect 1056 1491 1067 1537
rect 1113 1491 1124 1502
rect 2992 1501 3003 1547
rect 3196 1501 3207 1547
rect 3400 1501 3411 1547
rect 3604 1501 3615 1547
rect 3808 1501 3819 1547
rect 4012 1501 4023 1547
rect 260 -510 281 -499
rect 399 -510 420 -499
rect 1010 -540 1031 -529
rect 1149 -540 1170 -529
rect 306 -591 317 -545
rect 1056 -621 1067 -575
rect 3196 -611 3207 -565
rect 3400 -611 3411 -565
rect 3604 -611 3615 -565
rect 3808 -611 3819 -565
rect 4012 -611 4023 -565
rect 4752 -910 4766 4216
rect 4830 -910 4844 4216
rect 4908 -910 4922 4216
rect 4986 -910 5000 4216
rect 5064 -910 5078 4216
rect 5142 -910 5156 4216
rect 5220 -910 5234 4216
rect 5298 -910 5312 4216
rect 5376 -910 5390 4216
rect 5454 -910 5468 4216
rect 5532 -910 5546 4216
rect 5610 -910 5624 4216
rect 5688 -910 5702 4216
rect 5766 -910 5780 4216
rect 5844 -910 5858 4216
rect 5922 -910 5936 4216
rect 6000 -910 6014 4216
rect 6078 -910 6092 4216
rect 6156 -910 6170 4216
rect 6234 -910 6248 4216
rect 6312 -910 6326 4216
rect 6390 -910 6404 4216
rect 6468 -910 6482 4216
rect 6546 -910 6560 4216
rect 6624 -910 6638 4216
rect 6702 -910 6716 4216
rect 6780 -910 6794 4216
rect 6858 -910 6872 4216
rect 6936 -910 6950 4216
rect 7014 -910 7028 4216
rect 7092 -910 7106 4216
rect 7170 -910 7184 4216
rect 7248 -910 7262 4216
rect 7326 -910 7340 4216
rect 7404 -910 7418 4216
rect 7482 -910 7496 4216
rect 7560 -910 7574 4216
rect 7638 -910 7652 4216
rect 7716 -910 7730 4216
rect 7794 -910 7808 4216
rect 7872 -910 7886 4216
rect 7950 -910 7964 4216
rect 8028 -910 8042 4216
rect 8106 -910 8120 4216
rect 8184 -910 8198 4216
rect 8262 -910 8276 4216
rect 8340 -910 8354 4216
rect 8418 -910 8432 4216
rect 8496 -910 8510 4216
rect 8574 -910 8588 4216
rect 8652 -910 8666 4216
rect 8730 -910 8744 4216
rect 8808 -910 8822 4216
rect 8886 -910 8900 4216
rect 8964 -910 8978 4216
rect 9042 -910 9056 4216
rect 9120 -910 9134 4216
rect 9198 -910 9212 4216
rect 9276 -910 9290 4216
rect 9354 -910 9368 4216
rect 9432 -910 9446 4216
rect 9510 -910 9524 4216
rect 9588 -910 9602 4216
rect 9666 -910 9680 4216
rect 9744 -910 9758 4216
rect 9822 -910 9836 4216
rect 9900 -910 9914 4216
rect 9978 -910 9992 4216
rect -658 -2920 -644 -1354
rect -580 -2920 -566 -1354
rect -502 -2920 -488 -1354
rect -424 -2920 -410 -1354
rect -346 -2920 -332 -1354
rect -268 -2920 -254 -1354
rect -190 -2920 -176 -1354
rect -112 -2920 -98 -1354
rect -34 -2920 -20 -1354
rect 44 -2920 58 -1354
rect 122 -2920 136 -1354
rect 200 -2920 214 -1354
rect 278 -2920 292 -1354
rect 356 -2920 370 -1354
rect 434 -2920 448 -1354
rect 512 -2920 526 -1354
rect 590 -2920 604 -1354
rect 668 -2920 682 -1354
rect 746 -2920 760 -1354
rect 824 -2920 838 -1354
rect 902 -2920 916 -1354
rect 980 -2920 994 -1354
rect 1058 -2920 1072 -1354
rect 1136 -2920 1150 -1354
rect 1214 -2920 1228 -1354
rect 1292 -2920 1306 -1354
rect 1370 -2920 1384 -1354
rect 1448 -2920 1462 -1354
rect 1526 -2920 1540 -1354
rect 1604 -2920 1618 -1354
rect 1682 -2920 1696 -1354
rect 1760 -2920 1774 -1354
rect 1838 -2920 1852 -1354
rect 1916 -2920 1930 -1354
rect 1994 -2920 2008 -1354
rect 2072 -2920 2086 -1354
rect 2150 -2920 2164 -1354
rect 2228 -2920 2242 -1354
rect 2306 -2920 2320 -1354
rect 2384 -2920 2398 -1354
rect 2462 -2920 2476 -1354
rect 2540 -2920 2554 -1354
rect 2618 -2920 2632 -1354
rect 2696 -2920 2710 -1354
rect 2774 -2920 2788 -1354
rect 2852 -2920 2866 -1354
rect 2930 -2920 2944 -1354
rect 3008 -2920 3022 -1354
rect 3086 -2920 3100 -1354
rect 3164 -2920 3178 -1354
rect 3242 -2920 3256 -1354
rect 3320 -2920 3334 -1354
rect 3398 -2920 3412 -1354
rect 3476 -2920 3490 -1354
rect 3554 -2920 3568 -1354
rect 3632 -2920 3646 -1354
rect 3710 -2920 3724 -1354
rect 3788 -2920 3802 -1354
rect 3866 -2920 3880 -1354
rect 3944 -2920 3958 -1354
rect 4022 -2920 4036 -1354
rect 4100 -2920 4114 -1354
rect 4178 -2920 4192 -1354
rect 4256 -2920 4270 -1354
rect 4334 -2920 4348 -1354
rect 4412 -2920 4426 -1354
rect 4490 -2920 4504 -1354
rect 4568 -2920 4582 -1354
rect 4646 -2920 4660 -1354
rect 4724 -2920 4738 -1354
rect 4802 -2920 4816 -1354
rect 4880 -2920 4894 -1354
rect 4958 -2920 4972 -1354
rect 5036 -2920 5050 -1354
rect 5114 -2920 5128 -1354
rect 5192 -2920 5206 -1354
rect 5270 -2920 5284 -1354
rect 5348 -2920 5362 -1354
rect 5426 -2920 5440 -1354
rect 5504 -2920 5518 -1354
rect 5582 -2920 5596 -1354
rect 5660 -2920 5674 -1354
rect 5738 -2920 5752 -1354
rect 5816 -2920 5830 -1354
rect 5894 -2920 5908 -1354
rect 5972 -2920 5986 -1354
rect 6050 -2920 6064 -1354
rect 6128 -2920 6142 -1354
rect 6206 -2920 6220 -1354
rect 6284 -2920 6298 -1354
rect 6362 -2920 6376 -1354
rect 6440 -2920 6454 -1354
rect 6518 -2920 6532 -1354
rect 6596 -2920 6610 -1354
rect 6674 -2920 6688 -1354
rect 6752 -2920 6766 -1354
rect 6830 -2920 6844 -1354
rect 6908 -2920 6922 -1354
rect 6986 -2920 7000 -1354
rect 7064 -2920 7078 -1354
rect 7142 -2920 7156 -1354
rect 7220 -2920 7234 -1354
rect 7298 -2920 7312 -1354
rect 7376 -2920 7390 -1354
rect 7454 -2920 7468 -1354
rect 7532 -2920 7546 -1354
rect 7610 -2920 7624 -1354
rect 7688 -2920 7702 -1354
rect 7766 -2920 7780 -1354
rect 7844 -2920 7858 -1354
rect 7922 -2920 7936 -1354
rect 8000 -2920 8014 -1354
rect 8078 -2920 8092 -1354
rect 8156 -2920 8170 -1354
rect 8234 -2920 8248 -1354
rect 8312 -2920 8326 -1354
rect 8390 -2920 8404 -1354
rect 8468 -2920 8482 -1354
rect 8546 -2920 8560 -1354
rect 8624 -2920 8638 -1354
rect 8702 -2920 8716 -1354
rect 8780 -2920 8794 -1354
rect 8858 -2920 8872 -1354
rect 8936 -2920 8950 -1354
rect 9014 -2920 9028 -1354
rect 9092 -2920 9106 -1354
rect 9170 -2920 9184 -1354
rect 9248 -2920 9262 -1354
rect 9326 -2920 9340 -1354
rect 9404 -2920 9418 -1354
rect 9482 -2920 9496 -1354
rect 9560 -2920 9574 -1354
rect 9638 -2920 9652 -1354
rect 9716 -2920 9730 -1354
rect 9794 -2920 9808 -1354
rect 9872 -2920 9886 -1354
<< metal1 >>
rect -210 4180 3170 4370
rect 60 4060 90 4120
rect 150 4060 180 4120
rect 990 4060 1020 4120
rect 1090 4060 1110 4120
rect -170 2260 10 4040
rect 190 2890 210 3500
rect 280 2890 300 3500
rect 880 2890 900 3500
rect 960 2890 980 3500
rect 1160 2260 1340 4040
rect 1540 2630 1780 3500
rect 360 -70 380 1020
rect 460 -70 480 1020
rect 950 70 970 830
rect 1040 70 1060 830
rect 1120 -80 1140 990
rect 1210 -80 1230 990
rect 2320 -150 2530 610
rect 4090 -150 4330 620
rect -540 -340 -460 -300
rect -550 -450 -540 -340
rect -460 -450 -450 -340
rect -540 -480 -460 -450
rect -290 -530 -90 -220
rect -430 -620 -410 -560
rect -350 -620 -330 -560
rect 1820 -620 1860 -560
rect 1930 -620 1970 -560
rect 2130 -620 2170 -560
rect 2240 -620 2280 -560
rect 3010 -610 3070 -540
rect -700 -920 4350 -670
<< via1 >>
rect 90 4060 150 4120
rect 1020 4060 1090 4120
rect 210 2890 280 3500
rect 900 2890 960 3500
rect 380 -70 460 1020
rect 970 70 1040 830
rect 1140 -80 1210 990
rect -540 -450 -460 -340
rect -410 -620 -350 -560
rect 1860 -620 1930 -560
rect 2170 -620 2240 -560
<< metal2 >>
rect 40 4120 200 4400
rect 40 4060 90 4120
rect 150 4060 200 4120
rect 970 4120 1130 4360
rect 970 4060 1020 4120
rect 1090 4060 1130 4120
rect 40 4050 180 4060
rect 970 4050 1130 4060
rect 180 3500 310 3510
rect 180 2890 210 3500
rect 280 2890 310 3500
rect 180 1250 310 2890
rect 860 3500 980 3510
rect 860 2890 900 3500
rect 960 2890 980 3500
rect 860 1980 980 2890
rect 860 1850 1060 1980
rect 360 1020 610 1040
rect 360 -70 380 1020
rect 460 -70 490 1020
rect 590 -70 610 1020
rect 950 830 1060 1850
rect 950 70 970 830
rect 1040 70 1060 830
rect 950 40 1060 70
rect 1120 990 1340 1010
rect 360 -90 610 -70
rect 1120 -80 1140 990
rect 1210 -80 1250 990
rect 1330 -80 1340 990
rect 1120 -100 1340 -80
rect -550 -340 -330 -330
rect -550 -450 -540 -340
rect -460 -450 -330 -340
rect -550 -460 -330 -450
rect -430 -560 -330 -460
rect -430 -620 -410 -560
rect -350 -620 -330 -560
rect -430 -750 -330 -620
rect 1800 -560 2300 -540
rect 1800 -620 1860 -560
rect 1930 -620 2170 -560
rect 2240 -620 2300 -560
rect 1800 -640 2300 -620
rect 2000 -750 2100 -640
rect -430 -860 2100 -750
<< via2 >>
rect 490 -70 590 1020
rect 1250 -80 1330 990
<< metal3 >>
rect 480 -70 490 1020
rect 590 990 1340 1020
rect 590 -70 1250 990
rect 1240 -80 1250 -70
rect 1330 -80 1340 990
use mim_2p0fF_57EW3L  mim_2p0fF_57EW3L_0
timestamp 1691291836
transform 1 0 4820 0 1 6890
box -5240 -2120 5240 2120
use nmos_3p3_4JTTUB  nmos_3p3_4JTTUB_0
timestamp 1691291836
transform 1 0 2052 0 1 258
box -502 -1008 502 1008
use nmos_3p3_6FW5EE  nmos_3p3_6FW5EE_0
timestamp 1691270469
transform 1 0 3550 0 1 468
box -810 -1208 810 1208
use nmos_3p3_DTV5EE  nmos_3p3_DTV5EE_0
timestamp 1691270469
transform 1 0 1090 0 1 458
box -280 -1208 280 1208
use nmos_3p3_DTV5EE  nmos_3p3_DTV5EE_1
timestamp 1691270469
transform 1 0 340 0 1 488
box -280 -1208 280 1208
use nmos_3p3_VSY5LG  nmos_3p3_VSY5LG_0
timestamp 1691270469
transform 1 0 -380 0 1 -376
box -320 -374 320 374
use pmos_3p3_MAPLF9  pmos_3p3_MAPLF9_0
timestamp 1691436558
transform 1 0 4608 0 1 6888
box -5078 -2208 5078 2208
use pmos_3p3_TQ6DQ2  pmos_3p3_TQ6DQ2_0
timestamp 1691270469
transform 1 0 1050 0 1 3148
box -330 -1108 330 1108
use pmos_3p3_TQ6DQ2  pmos_3p3_TQ6DQ2_1
timestamp 1691270469
transform 1 0 120 0 1 3148
box -330 -1108 330 1108
use pmos_3p3_Z53MQA  pmos_3p3_Z53MQA_0
timestamp 1691270469
transform 1 0 2290 0 1 3038
box -750 -1208 750 1208
use rm1_8TUMYM  rm1_8TUMYM_0
timestamp 1691437249
transform 1 0 7349 0 1 1653
box -2629 -2563 2643 2563
use rm1_G26CKV  rm1_G26CKV_0
timestamp 1691437249
transform 1 0 4591 0 1 -3917
box -5281 -2563 5295 2563
<< end >>
