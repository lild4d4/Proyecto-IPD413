** Miller OTA Parameters **
.param otag=10
