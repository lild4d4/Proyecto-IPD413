** Bandgap Reference Parameters **

.param bgrv=1.2
